67.2987u
19.4695uupdate 222sp
fdfdfd.param vin='0.1'
